module try1
#(
parameter param1 = 3, parameter param2 = 4 
)
(
input [4:0] var1,
input [0:3] var2
);


endmodule
